//ejemplo de uso del módulo bluetooth HC06 como receptor
//adaptado a reloj de 25 MHz
///////////////////////////////////////////////////
module top(
    input clk,             //25MHz
    input reset,
    input rx,
    output reg [7:0] leds,
    output reg IO1, // Ahora son regs para poder resetearlos
    output reg IO2, // Ahora son regs para poder resetearlos
    output reg IO3, // Ahora son regs para poder resetearlos
    output reg IO4, // Ahora son regs para poder resetearlos
    output reg PWM,
    output reg PWM2
    
);

//fsm states
reg [1:0] presentstate, nextstate;
parameter EDO_1 = 2'b00;
parameter EDO_2 = 2'b10;

//señales
reg control=0;
reg done=0;
reg [8:0] tmp = 9'b000000000;

//contadores
reg [3:0] i = 4'b0000;
reg [8:0] c = 9'b111111111;    // <-- ajustado para 25 MHz
reg delay = 0;
reg [1:0] c2 = 2'b11;
reg capture = 0;
reg [19:0] cnt= 0;
always @(posedge clk) cnt <= cnt+1;


// ---------------------------------------------
// Retardo para reloj 25MHz
// c < 434  → 434 * 40ns ≈ 17.36us
// triple → ~52us
// doble → ~104us = 9600 baudios
// ---------------------------------------------
always @(posedge clk)
begin
    if(c < 9'd434)
        c = c + 1;
    else begin
        c = 0;
        delay = ~delay;
    end
end

// contador c2
always @(posedge delay)
begin
    if (c2 > 1)
        c2 = 0;
    else
        c2 = c2 + 1;
end

// captura
always @(c2)
begin
    if (c2 == 1)
        capture = 1;
    else
        capture = 0;
end

// FSM actualiza
always @(posedge capture or posedge reset)
begin
    if (reset)
        presentstate <= EDO_1;
    else
        presentstate <= nextstate;
end

// FSM lógica
always @(*)
begin
    case(presentstate)
    EDO_1:
        if(rx==1 && done==0) begin
            control = 0;
            nextstate = EDO_1;
        end 
        else if(rx==0 && done==0) begin
            control = 1;
            nextstate = EDO_2;
        end 
        else begin
            control = 0;
            nextstate = EDO_1;
        end

    EDO_2:
        if(done==0) begin
            control = 1;
            nextstate = EDO_2;
        end
        else begin
            control = 0;
            nextstate = EDO_1;
        end

    default: nextstate = EDO_1;
    endcase
end

// recepción de bits
always @(posedge capture)
begin
    if (control==1 && done==0)
        tmp <= {rx, tmp[8:1]};
end

// contador de bits
always @(posedge capture)
begin
    if (control) begin
        if(i >= 9) begin
            i = 0;
            done = 1;
            leds <= tmp[8:1];
        end
        else begin
            i = i + 1;
            done = 0;
        end
    end 
    else done = 0;
end

// --- LÓGICA DE CONTROL DE MOTORES Y PWM (Corregida) ---

reg [7:0] duty = 0;
reg [7:0] duty2 = 0;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        // Asegurar que todo se detenga al resetear
        IO1 <= 0;
        IO2 <= 0;
        IO3 <= 0;
        IO4 <= 0;
        duty <= 0;
        duty2 <= 0;
    end
    else begin
        case (leds)
            // 'A' -> Adelante (Velocidad media/alta)
            "A": begin
                IO1 <= 1; // Motor Derecho (M1) Forward
                IO2 <= 0;
                IO3 <= 1; // Motor Izquierdo (M2) Forward
                IO4 <= 0;
                duty <= 8'd90;  // PWM Motor Derecho
                duty2 <= 8'd90; // PWM Motor Izquierdo
            end
            
            // 'C' -> Detener (Stop/Frenado)
            "C": begin
                IO1 <= 0;
                IO2 <= 0;
                IO3 <= 0;
                IO4 <= 0;
                duty <= 8'd0;
                duty2 <= 8'd0;
            end
            
            // 'B' -> Retroceso (Velocidad media/alta)
            "B": begin
                IO1 <= 0; // Motor Derecho Reverse
                IO2 <= 1;
                IO3 <= 0; // Motor Izquierdo Reverse
                IO4 <= 1;
                duty <= 8'd90;
                duty2 <= 8'd90;
            end

            // 'F' -> Superior Derecha (Forward-Right Diagonal)
            "F": begin
                IO1 <= 1; // Motor Derecho Forward
                IO2 <= 0;
                IO3 <= 1; // Motor Izquierdo Forward
                IO4 <= 0;
                duty <= 8'd90;   // M1 (Derecho) Lento
                duty2 <= 8'd60; // M2 (Izquierdo) Rápido -> Gira a la derecha
            end
            
            // 'D' -> Girar a la Derecha (Pivot Derecha)
            "D": begin
                IO1 <= 0; // Motor Derecho (M1) Detenido (o Lento)
                IO2 <= 0;
                IO3 <= 1; // Motor Izquierdo (M2) Forward
                IO4 <= 0;
                duty <= 8'd90;   // Velocidad para M1 (aunque IOs lo detienen)
                duty2 <= 8'd155; // Velocidad para M2
            end

            // === NUEVA LÓGICA ===
            
            // 'G' -> Superior Izquierda (Forward-Left Diagonal)
            "E": begin
                IO1 <= 1; // Motor Derecho (M1) Forward
                IO2 <= 0;
                IO3 <= 1; // Motor Izquierdo (M2) Forward
                IO4 <= 0;
                duty <= 8'd90; // M1 (Derecho) Rápido -> Gira a la izquierda
                duty2 <= 8'd60;  // M2 (Izquierdo) Lento
            end
            
            // 'I' -> Girar Izquierda (Spin/Pivot Izquierda)
            "G": begin
                IO1 <= 1; // Motor Derecho (M1) Forward
                IO2 <= 0;
                IO3 <= 0; // Motor Izquierdo (M2) Reverse
                IO4 <= 1;
                duty <= 8'd90;  // M1 (Derecho)
                duty2 <= 8'd90; // M2 (Izquierdo) - Misma velocidad para giro cerrado
            end
            
            default: begin
                // Mantener el estado
            end
        endcase
    end
end

// Generación de la señal PWM 1
// PWM es 'alto' mientras el contador 'cnt' esté por debajo de 'duty'
always @(posedge clk)
    PWM <= (cnt[18:11] < duty);

// Generación de la señal PWM 2
always @(posedge clk)
    PWM2 <= (cnt[18:11] < duty2);

endmodule
